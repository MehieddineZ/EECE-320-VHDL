Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity mux8to1_TB is
end mux8to1_TB;
Architecture mux8to1_TB_arch of  mux8to1_TB is 

component mux8to1 is 
port(
	S :  IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	I0,I1,I2,I3,I4,I5,I6,I7,G : IN STD_LOGIC;
	F: OUT STD_LOGIC

);
end component;
signal I0,I1,I2,I3,I4,I5,I6,I7,G,F : STD_LOGIC := '0';
signal S: STD_LOGIC_VECTOR(2 downto 0);
begin
      UUT: mux8to1 Port Map (S=>S,I0=>I0 , I1=>I1 , I2=>I2 ,I3=>I3,I4=>I4 ,I5=>I5 ,I6=>I6,I7=>I7,G=>G,F=>F);
         PROCESS
		BEGIN
			

		G<='1';
		S<="000";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
			
		S<="001";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="010";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="011";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;

	S<="100";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="101";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="110";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="111";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	G<='0';
		S<="000";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
			
		S<="001";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="010";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="011";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;

	S<="100";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="101";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="110";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
	S<="111";
			I0<='1'; 
			wait for 10ns;
			I0<='0';
			wait for 10ns;
			I1<='1';
			wait for 10ns;
			I1<='0';
			wait for 10ns;
			I2<='1';
			wait for 10ns;
			I2<='0';
			wait for 10ns;
			I3<='1' ;
			wait for 10ns;
			I3<='0';
			wait for 10ns;
			I4<='1';
			wait for 10ns;
			I4<='0';
			wait for 10ns;
			I5<='1' ;
			wait for 10ns;
			I5<='0' ;
			wait for 10ns;
			I6<='1' ;
			wait for 10ns;
			I6<='0' ;
			wait for 10ns;
			I7<='1' ;
			wait for 10ns;
			I7<='0' ;
wait;
end PROCESS;
end mux8to1_TB_arch;
			
			
			
			
			
			
			